`timescale 1ns/100ps
module rom(clk, data, addr);
output [23:0] data;
input [8:0] addr;
input clk;

reg [23:0] data;
reg [23:0] romdata;

always @(posedge clk) begin
	data <= romdata;
end

// 22 bit FP
always @(addr) begin
	case (addr)
		0: romdata = 663;
		1: romdata = 215;
		2: romdata = 194;
		3: romdata = 130;
		4: romdata = 27;
		5: romdata = -106;
		6: romdata = -252;
		7: romdata = -389;
		8: romdata = -492;
		9: romdata = -539;
		10: romdata = -514;
		11: romdata = -412;
		12: romdata = -238;
		13: romdata = -11;
		14: romdata = 239;
		15: romdata = 473;
		16: romdata = 651;
		17: romdata = 738;
		18: romdata = 707;
		19: romdata = 551;
		20: romdata = 280;
		21: romdata = -75;
		22: romdata = -464;
		23: romdata = -827;
		24: romdata = -1101;
		25: romdata = -1233;
		26: romdata = -1183;
		27: romdata = -941;
		28: romdata = -524;
		29: romdata = 17;
		30: romdata = 608;
		31: romdata = 1159;
		32: romdata = 1577;
		33: romdata = 1779;
		34: romdata = 1714;
		35: romdata = 1365;
		36: romdata = 761;
		37: romdata = -24;
		38: romdata = -880;
		39: romdata = -1677;
		40: romdata = -2280;
		41: romdata = -2575;
		42: romdata = -2487;
		43: romdata = -1994;
		44: romdata = -1142;
		45: romdata = -34;
		46: romdata = 1173;
		47: romdata = 2295;
		48: romdata = 3145;
		49: romdata = 3565;
		50: romdata = 3451;
		51: romdata = 2779;
		52: romdata = 1610;
		53: romdata = 91;
		54: romdata = -1564;
		55: romdata = -3102;
		56: romdata = -4268;
		57: romdata = -4849;
		58: romdata = -4706;
		59: romdata = -3807;
		60: romdata = -2238;
		61: romdata = -198;
		62: romdata = 2025;
		63: romdata = 4090;
		64: romdata = 5658;
		65: romdata = 6445;
		66: romdata = 6270;
		67: romdata = 5092;
		68: romdata = 3026;
		69: romdata = 338;
		70: romdata = -2590;
		71: romdata = -5312;
		72: romdata = -7382;
		73: romdata = -8429;
		74: romdata = -8218;
		75: romdata = -6698;
		76: romdata = -4023;
		77: romdata = -539;
		78: romdata = 3259;
		79: romdata = 6789;
		80: romdata = 9479;
		81: romdata = 10850;
		82: romdata = 10602;
		83: romdata = 8671;
		84: romdata = 5256;
		85: romdata = 803;
		86: romdata = -4052;
		87: romdata = -8568;
		88: romdata = -12015;
		89: romdata = -13785;
		90: romdata = -13498;
		91: romdata = -11076;
		92: romdata = -6772;
		93: romdata = -1153;
		94: romdata = 4978;
		95: romdata = 10685;
		96: romdata = 15049;
		97: romdata = 17306;
		98: romdata = 16981;
		99: romdata = 13977;
		100: romdata = 8615;
		101: romdata = 1601;
		102: romdata = -6056;
		103: romdata = -13191;
		104: romdata = -18656;
		105: romdata = -21504;
		106: romdata = -21143;
		107: romdata = -17455;
		108: romdata = -10839;
		109: romdata = -2171;
		110: romdata = 7300;
		111: romdata = 16135;
		112: romdata = 22917;
		113: romdata = 26475;
		114: romdata = 26084;
		115: romdata = 21598;
		116: romdata = 13506;
		117: romdata = 2886;
		118: romdata = -8731;
		119: romdata = -19580;
		120: romdata = -27927;
		121: romdata = -32338;
		122: romdata = -31925;
		123: romdata = -26511;
		124: romdata = -16689;
		125: romdata = -3774;
		126: romdata = 10371;
		127: romdata = 23599;
		128: romdata = 33799;
		129: romdata = 39229;
		130: romdata = 38809;
		131: romdata = 32319;
		132: romdata = 20477;
		133: romdata = 4870;
		134: romdata = -12248;
		135: romdata = -28279;
		136: romdata = -40672;
		137: romdata = -47320;
		138: romdata = -46912;
		139: romdata = -39179;
		140: romdata = -24977;
		141: romdata = -6216;
		142: romdata = 14395;
		143: romdata = 33731;
		144: romdata = 48720;
		145: romdata = 56823;
		146: romdata = 56457;
		147: romdata = 47285;
		148: romdata = 30328;
		149: romdata = 7866;
		150: romdata = -16858;
		151: romdata = -40099;
		152: romdata = -58169;
		153: romdata = -68018;
		154: romdata = -67735;
		155: romdata = -56898;
		156: romdata = -36712;
		157: romdata = -9889;
		158: romdata = 19700;
		159: romdata = 47577;
		160: romdata = 69326;
		161: romdata = 81284;
		162: romdata = 81141;
		163: romdata = 68369;
		164: romdata = 44375;
		165: romdata = 12380;
		166: romdata = -23007;
		167: romdata = -56436;
		168: romdata = -82618;
		169: romdata = -97149;
		170: romdata = -97233;
		171: romdata = -82192;
		172: romdata = -53667;
		173: romdata = -15470;
		174: romdata = 26906;
		175: romdata = 67068;
		176: romdata = 98667;
		177: romdata = 116388;
		178: romdata = 116827;
		179: romdata = 99100;
		180: romdata = 65105;
		181: romdata = 19357;
		182: romdata = -31593;
		183: romdata = -80070;
		184: romdata = -118419;
		185: romdata = -140185;
		186: romdata = -141177;
		187: romdata = -120220;
		188: romdata = -79491;
		189: romdata = -24341;
		190: romdata = 37376;
		191: romdata = 96392;
		192: romdata = 143393;
		193: romdata = 170450;
		194: romdata = 172322;
		195: romdata = 147400;
		196: romdata = 98147;
		197: romdata = 30924;
		198: romdata = -44780;
		199: romdata = -117648;
		200: romdata = -176185;
		201: romdata = -210477;
		202: romdata = -213812;
		203: romdata = -183886;
		204: romdata = -123414;
		205: romdata = -39997;
		206: romdata = 54762;
		207: romdata = 146804;
		208: romdata = 221623;
		209: romdata = 266471;
		210: romdata = 272414;
		211: romdata = 235949;
		212: romdata = 159885;
		213: romdata = 53333;
		214: romdata = -69263;
		215: romdata = -189961;
		216: romdata = -289806;
		217: romdata = -351634;
		218: romdata = -362805;
		219: romdata = -317461;
		220: romdata = -217928;
		221: romdata = -75021;
		222: romdata = 92878;
		223: romdata = 261932;
		224: romdata = 405905;
		225: romdata = 499834;
		226: romdata = 523805;
		227: romdata = 466342;
		228: romdata = 326904;
		229: romdata = 117086;
		230: romdata = -139721;
		231: romdata = -410270;
		232: romdata = -654846;
		233: romdata = -831751;
		234: romdata = -902362;
		235: romdata = -836171;
		236: romdata = -615143;
		237: romdata = -236839;
		238: romdata = 284164;
		239: romdata = 916784;
		240: romdata = 1615898;
		241: romdata = 2326541;
		242: romdata = 2989376;
		243: romdata = 3546834;
		244: romdata = 3949221;
		245: romdata = 4160060;
		246: romdata = 4160060;
		247: romdata = 3949221;
		248: romdata = 3546834;
		249: romdata = 2989376;
		250: romdata = 2326541;
		251: romdata = 1615898;
		252: romdata = 916784;
		253: romdata = 284164;
		254: romdata = -236839;
		255: romdata = -615143;
		256: romdata = -836171;
		257: romdata = -902362;
		258: romdata = -831751;
		259: romdata = -654846;
		260: romdata = -410270;
		261: romdata = -139721;
		262: romdata = 117086;
		263: romdata = 326904;
		264: romdata = 466342;
		265: romdata = 523805;
		266: romdata = 499834;
		267: romdata = 405905;
		268: romdata = 261932;
		269: romdata = 92878;
		270: romdata = -75021;
		271: romdata = -217928;
		272: romdata = -317461;
		273: romdata = -362805;
		274: romdata = -351634;
		275: romdata = -289806;
		276: romdata = -189961;
		277: romdata = -69263;
		278: romdata = 53333;
		279: romdata = 159885;
		280: romdata = 235949;
		281: romdata = 272414;
		282: romdata = 266471;
		283: romdata = 221623;
		284: romdata = 146804;
		285: romdata = 54762;
		286: romdata = -39997;
		287: romdata = -123414;
		288: romdata = -183886;
		289: romdata = -213812;
		290: romdata = -210477;
		291: romdata = -176185;
		292: romdata = -117648;
		293: romdata = -44780;
		294: romdata = 30924;
		295: romdata = 98147;
		296: romdata = 147400;
		297: romdata = 172322;
		298: romdata = 170450;
		299: romdata = 143393;
		300: romdata = 96392;
		301: romdata = 37376;
		302: romdata = -24341;
		303: romdata = -79491;
		304: romdata = -120220;
		305: romdata = -141177;
		306: romdata = -140185;
		307: romdata = -118419;
		308: romdata = -80070;
		309: romdata = -31593;
		310: romdata = 19357;
		311: romdata = 65105;
		312: romdata = 99100;
		313: romdata = 116827;
		314: romdata = 116388;
		315: romdata = 98667;
		316: romdata = 67068;
		317: romdata = 26906;
		318: romdata = -15470;
		319: romdata = -53667;
		320: romdata = -82192;
		321: romdata = -97233;
		322: romdata = -97149;
		323: romdata = -82618;
		324: romdata = -56436;
		325: romdata = -23007;
		326: romdata = 12380;
		327: romdata = 44375;
		328: romdata = 68369;
		329: romdata = 81141;
		330: romdata = 81284;
		331: romdata = 69326;
		332: romdata = 47577;
		333: romdata = 19700;
		334: romdata = -9889;
		335: romdata = -36712;
		336: romdata = -56898;
		337: romdata = -67735;
		338: romdata = -68018;
		339: romdata = -58169;
		340: romdata = -40099;
		341: romdata = -16858;
		342: romdata = 7866;
		343: romdata = 30328;
		344: romdata = 47285;
		345: romdata = 56457;
		346: romdata = 56823;
		347: romdata = 48720;
		348: romdata = 33731;
		349: romdata = 14395;
		350: romdata = -6216;
		351: romdata = -24977;
		352: romdata = -39179;
		353: romdata = -46912;
		354: romdata = -47320;
		355: romdata = -40672;
		356: romdata = -28279;
		357: romdata = -12248;
		358: romdata = 4870;
		359: romdata = 20477;
		360: romdata = 32319;
		361: romdata = 38809;
		362: romdata = 39229;
		363: romdata = 33799;
		364: romdata = 23599;
		365: romdata = 10371;
		366: romdata = -3774;
		367: romdata = -16689;
		368: romdata = -26511;
		369: romdata = -31925;
		370: romdata = -32338;
		371: romdata = -27927;
		372: romdata = -19580;
		373: romdata = -8731;
		374: romdata = 2886;
		375: romdata = 13506;
		376: romdata = 21598;
		377: romdata = 26084;
		378: romdata = 26475;
		379: romdata = 22917;
		380: romdata = 16135;
		381: romdata = 7300;
		382: romdata = -2171;
		383: romdata = -10839;
		384: romdata = -17455;
		385: romdata = -21143;
		386: romdata = -21504;
		387: romdata = -18656;
		388: romdata = -13191;
		389: romdata = -6056;
		390: romdata = 1601;
		391: romdata = 8615;
		392: romdata = 13977;
		393: romdata = 16981;
		394: romdata = 17306;
		395: romdata = 15049;
		396: romdata = 10685;
		397: romdata = 4978;
		398: romdata = -1153;
		399: romdata = -6772;
		400: romdata = -11076;
		401: romdata = -13498;
		402: romdata = -13785;
		403: romdata = -12015;
		404: romdata = -8568;
		405: romdata = -4052;
		406: romdata = 803;
		407: romdata = 5256;
		408: romdata = 8671;
		409: romdata = 10602;
		410: romdata = 10850;
		411: romdata = 9479;
		412: romdata = 6789;
		413: romdata = 3259;
		414: romdata = -539;
		415: romdata = -4023;
		416: romdata = -6698;
		417: romdata = -8218;
		418: romdata = -8429;
		419: romdata = -7382;
		420: romdata = -5312;
		421: romdata = -2590;
		422: romdata = 338;
		423: romdata = 3026;
		424: romdata = 5092;
		425: romdata = 6270;
		426: romdata = 6445;
		427: romdata = 5658;
		428: romdata = 4090;
		429: romdata = 2025;
		430: romdata = -198;
		431: romdata = -2238;
		432: romdata = -3807;
		433: romdata = -4706;
		434: romdata = -4849;
		435: romdata = -4268;
		436: romdata = -3102;
		437: romdata = -1564;
		438: romdata = 91;
		439: romdata = 1610;
		440: romdata = 2779;
		441: romdata = 3451;
		442: romdata = 3565;
		443: romdata = 3145;
		444: romdata = 2295;
		445: romdata = 1173;
		446: romdata = -34;
		447: romdata = -1142;
		448: romdata = -1994;
		449: romdata = -2487;
		450: romdata = -2575;
		451: romdata = -2280;
		452: romdata = -1677;
		453: romdata = -880;
		454: romdata = -24;
		455: romdata = 761;
		456: romdata = 1365;
		457: romdata = 1714;
		458: romdata = 1779;
		459: romdata = 1577;
		460: romdata = 1159;
		461: romdata = 608;
		462: romdata = 17;
		463: romdata = -524;
		464: romdata = -941;
		465: romdata = -1183;
		466: romdata = -1233;
		467: romdata = -1101;
		468: romdata = -827;
		469: romdata = -464;
		470: romdata = -75;
		471: romdata = 280;
		472: romdata = 551;
		473: romdata = 707;
		474: romdata = 738;
		475: romdata = 651;
		476: romdata = 473;
		477: romdata = 239;
		478: romdata = -11;
		479: romdata = -238;
		480: romdata = -412;
		481: romdata = -514;
		482: romdata = -539;
		483: romdata = -492;
		484: romdata = -389;
		485: romdata = -252;
		486: romdata = -106;
		487: romdata = 27;
		488: romdata = 130;
		489: romdata = 194;
		490: romdata = 215;
		491: romdata = 663;
		default: romdata = 0;
	endcase
end

endmodule